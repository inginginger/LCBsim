module answers(
input clk80MHz,
input rst,
input addr,
output reg[7:0] data);

reg [7:0] cnt;

always@(posedge clk80MHz or negedge rst)
begin
	if(~rst) begin
		data <= 7'd0;
		cnt <= 8'd0;
	end
	else begin
		case(addr)
			0 : data <= cnt ;
			1 : data <= 7'd10;
			2 : data <= 7'd20;
			3 : data <= 7'd30;
			4 : data <= 7'd40;
			5 : data <= 7'd50;
			6 : data <= 7'd60;
			7 : data <= 7'd70;
			8 : data <= 7'd80;
			9 : data <= 7'd90;
			10 : data <= 7'd100;
			11 : data <= 7'd110;
			12 : data <= 7'd120;
			13 : data <= 7'd130;
			14 : data <= 7'd140;
			15 : data <= 7'd150;
			16 : data <= 7'd160;
			17 : data <= 7'd170;
			18 : data <= 7'd180;
			19 : begin
				data <= 7'd190;
				cnt <= cnt + 1;
				/*if(cnt == 8'd255)
					cnt <= 8'd0;*/
			end
		endcase
	end
end
endmodule